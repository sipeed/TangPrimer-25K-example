/*LED流水灯以及拨码开关真值显示模块*/
module driver_Led(
    input           i_clk               ,
    input           i_rst               ,
    input   [3:0]   i_switch            ,
    output  [7:0]   o_led
);
/***************reg*******************/
reg         [27:0]  r_cnt       = 0             ;
reg         [7:0]   r_streamLed = 8'b11111110   ;//输出流水灯寄存器
reg         [7:0]   w_tabelLed  = 8'b11111111   ;//输出拨码开关真值表寄存器
/***************assign****************/
assign      o_led = i_switch[3] ? w_tabelLed : r_streamLed;//当拨码开关的最高位(最左边)为高时，显示流水灯，否则显示低三位(右三个)拨码开关的真值表
/***************always****************/
//——————<w_tabelLed>—————————————//
always @(posedge i_clk or posedge i_rst)
begin
    if(i_rst)
        w_tabelLed  <= 8'b11111111;
    else
        case(i_switch[2:0])
            3'b111  : w_tabelLed <= 8'b11111111;
            3'b110  : w_tabelLed <= 8'b11111110;
            3'b101  : w_tabelLed <= 8'b11111101;
            3'b100  : w_tabelLed <= 8'b11111011;
            3'b011  : w_tabelLed <= 8'b11110111;
            3'b010  : w_tabelLed <= 8'b11101111;
            3'b001  : w_tabelLed <= 8'b11011111;
            3'b000  : w_tabelLed <= 8'b10111111;
            default : w_tabelLed <= 8'b11111111;
        endcase
end
//——————<r_cnt>—————————————//
always @(posedge i_clk or posedge i_rst)
begin
    if(i_rst)
        r_cnt <= 0;
    else if(r_cnt == 'd50_000_000)
        r_cnt <= 0;
    else
        r_cnt <= r_cnt + 1;
end
//——————<r_streamLed>—————————————//
always @(posedge i_clk or posedge i_rst)
begin
    if(i_rst)
        r_streamLed <= 8'b11111110;
    else if(r_cnt == 'd50_000_000)
        r_streamLed <= {r_streamLed[6:0],r_streamLed[7]};
    else
        r_streamLed <= r_streamLed;
end
endmodule
