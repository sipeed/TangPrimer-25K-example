//Copyright (C)2014-2023 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.9 Beta-5
//Part Number: GW5A-LV25MG121NES
//Device: GW5A-25
//Device Version: A
//Created Time: Sun Oct 29 21:03:01 2023

module Gowin_pROM (dout, clk, oce, ce, reset, ad);

output [31:0] dout;
input clk;
input oce;
input ce;
input reset;
input [10:0] ad;

wire [23:0] prom_inst_0_dout_w;
wire [23:0] prom_inst_1_dout_w;
wire [23:0] prom_inst_2_dout_w;
wire [23:0] prom_inst_3_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[23:0],dout[7:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 8;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'hBBBBBBBBBBBBBABBFECC00000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_01 = 256'h000000000000000000000000000000000000000000B3FDBBBBBBBBBBBBBBBBBB;
defparam prom_inst_0.INIT_RAM_02 = 256'hBBBBBBBBBBBABBFECD0000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000B3FDBBBBBBBBBBBBBBBBBBBB;
defparam prom_inst_0.INIT_RAM_04 = 256'hBBBBBBBBBABBFECC000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_05 = 256'h00000000000000000000000000000000000000B3FEBBBBBBBBBBBBBBBBBBBBBB;
defparam prom_inst_0.INIT_RAM_06 = 256'hDBDBDBDBDCFECD00000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_07 = 256'h000000000000000000000000000000000000B3FEBBBABBDBDBDBDBDBDBDBDBDB;
defparam prom_inst_0.INIT_RAM_08 = 256'hBBBBBBBBDBCD0000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_09 = 256'h0000000000000000000000000000000000B3FEBBBBBBBBBBBABBBBBBBBBBBBBB;
defparam prom_inst_0.INIT_RAM_0A = 256'h6363636342000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_0B = 256'h00000000000000000000000000000000B3FDBBBBBBFDAC006363636363636363;
defparam prom_inst_0.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_0D = 256'h000000000000000000000000000000B3FDBBBBBBBBFD6B000000000000000000;
defparam prom_inst_0.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_0F = 256'h0000000000000000000000000000B3FDBBBBBBBBBBFD8B000000000000000000;
defparam prom_inst_0.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_11 = 256'h00000000000000000000000000B3FEBBBBBBBBBBBBFD8B000000000000000000;
defparam prom_inst_0.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_13 = 256'h000000000000000000000000D4FEBBBBBBBBBBBBBBFD8B000000000000000000;
defparam prom_inst_0.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_15 = 256'h000000000000000000000000ACFDDBBABBBBBBBBBBFD8B000000000000000000;
defparam prom_inst_0.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_17 = 256'h000000000000000000000000008BFDDBBABBBBBBBBFD8B000000000000000000;
defparam prom_inst_0.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_19 = 256'h00000000000000000000000000008AFDDBBBBBBBBBFD8B000000000000000000;
defparam prom_inst_0.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_1B = 256'h0000000000000000000000000000008BFDDBBBBBBBFD6A000000000000000000;
defparam prom_inst_0.INIT_RAM_1C = 256'h8B6B6B6B8B8B6B6B6B8B8B6B8B8C630000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_1D = 256'h000000000000000000000000000000008BFDDBBBBBDC514A6B8B8B8B6B6B6B8B;
defparam prom_inst_0.INIT_RAM_1E = 256'hFDFDFDFDFDFDFDFDFDFDFDFDFDFF080000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_1F = 256'h00000000000000000000000000000000008BFDDBBBBADCFEFDFDFDFDFDFDFDFD;
defparam prom_inst_0.INIT_RAM_20 = 256'hBBBBBBBBBBBBBBBBBBBBBBBBBBFCE70000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_21 = 256'h000000000000000000000000000000000000ABFDDBBABBBBBBBBBBBBBBBBBBBB;
defparam prom_inst_0.INIT_RAM_22 = 256'hBBBBBBBBBBBBBBBBBBBBBBBBBBFCE70000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_23 = 256'h00000000000000000000000000000000000000ABFDDBBBBBBBBBBBBBBBBBBBBB;
defparam prom_inst_0.INIT_RAM_24 = 256'hBBBBBBBBBBBBBBBBBBBBBBBBBBFCE70000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000ACFEDBBABBBBBBBBBBBBBBBB;
defparam prom_inst_0.INIT_RAM_26 = 256'hBBBBBBBBBBBBBBBBBBBBBBBBBBFCE70000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_27 = 256'h000000000000000000000000000000000000000000ACFDDBBABBBBBBBBBBBBBB;
defparam prom_inst_0.INIT_RAM_28 = 256'hBBBBBBBBBBBBBBBBBBBBBBBBBBFCE70000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_29 = 256'h00000000000000000000000000000000000000000000ACFEDBBABBBBBBBBBBBB;
defparam prom_inst_0.INIT_RAM_2A = 256'hBBBBBBBBBBBBBBBBBBBBBBBBBBFCE70000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000ACFEDBBABBBBBBBBBB;
defparam prom_inst_0.INIT_RAM_2C = 256'hFDFDFDFDFDFDFDFDFDFDFDFDFDFE070000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_2D = 256'h000000000000000000000000000000000000000000000000ACFEFDFDFDFDFDFD;
defparam prom_inst_0.INIT_RAM_2E = 256'h72727272727272727272727292B3A40000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_2F = 256'h000000000000000000000000000000000000000000000000008BB37272727272;
defparam prom_inst_0.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000042;
defparam prom_inst_0.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_36 = 256'h000000000000000000000000000000000000000000000000000000000000004A;
defparam prom_inst_0.INIT_RAM_37 = 256'hC600000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000018;
defparam prom_inst_0.INIT_RAM_39 = 256'h9300000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3A = 256'h000000000000000000000000000000000000000000000000000000000000EEBB;
defparam prom_inst_0.INIT_RAM_3B = 256'hBB6B000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000EFBBBB;
defparam prom_inst_0.INIT_RAM_3D = 256'hBBBB8B0000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000424A17BBBBBB;
defparam prom_inst_0.INIT_RAM_3F = 256'hBBBBBBD608210000000000000000000000000000000000000000000000000000;

pROM prom_inst_1 (
    .DO({prom_inst_1_dout_w[23:0],dout[15:8]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_1.READ_MODE = 1'b0;
defparam prom_inst_1.BIT_WIDTH = 8;
defparam prom_inst_1.RESET_MODE = "SYNC";
defparam prom_inst_1.INIT_RAM_00 = 256'h7F7F7F7F7F7F7F7F7F654C505454545454545454545454545454545454545454;
defparam prom_inst_1.INIT_RAM_01 = 256'h54545454545454545454545454545454545454504C6E7F7F7F7F7F7F7F7F7F7F;
defparam prom_inst_1.INIT_RAM_02 = 256'h7F7F7F7F7F7F7F7F655054545454545454545454545454545454545454545454;
defparam prom_inst_1.INIT_RAM_03 = 256'h545454545454545454545454545454545454504C6E7F7F7F7F7F7F7F7F7F7F7F;
defparam prom_inst_1.INIT_RAM_04 = 256'h7F7F7F7F7F7F7F65505054545454545454545454545454545454545454545454;
defparam prom_inst_1.INIT_RAM_05 = 256'h5454545454545454545454545454545454504C6E7F7F7F7F7F7F7F7F7F7F7F7F;
defparam prom_inst_1.INIT_RAM_06 = 256'h7F7F7F7F7F7F6550545454545454545454545454545454545454545454545454;
defparam prom_inst_1.INIT_RAM_07 = 256'h54545454545454545454545454545454504C6E7F7F7F7F7F7F7F7F7F7F7F7F7F;
defparam prom_inst_1.INIT_RAM_08 = 256'h7B7B7B7F7F655050545454545454545454545454545454545454545454545454;
defparam prom_inst_1.INIT_RAM_09 = 256'h545454545454545454545454545454504C6E7F7F7F7F7F7B7B7B7B7B7B7B7B7B;
defparam prom_inst_1.INIT_RAM_0A = 256'h5454545450505454545454545454545454545454545454545454545454545454;
defparam prom_inst_1.INIT_RAM_0B = 256'h5454545454545454545454545454504C6E7F7F7F7F7F61505454545454545454;
defparam prom_inst_1.INIT_RAM_0C = 256'h5050505054545454545454545454545454545454545454545454545454545454;
defparam prom_inst_1.INIT_RAM_0D = 256'h54545454545454545454545454504C6E7F7F7F7F7F7F614C5450505050505050;
defparam prom_inst_1.INIT_RAM_0E = 256'h5454545454545454545454545454545454545454545454545454545454545454;
defparam prom_inst_1.INIT_RAM_0F = 256'h545454545454545454545454504C6E7F7F7F7F7F7F7F61505454545454545454;
defparam prom_inst_1.INIT_RAM_10 = 256'h5454545454545454545454545454545454545454545454545454545454545454;
defparam prom_inst_1.INIT_RAM_11 = 256'h5454545454545454545454544C6E7F7F7F7F7F7F7F7F61505454545454545454;
defparam prom_inst_1.INIT_RAM_12 = 256'h5454545454545454545454545454545454545454545454545454545454545454;
defparam prom_inst_1.INIT_RAM_13 = 256'h5454545454545454545454506E7F7F7F7F7F7F7F7F7F61505454545454545454;
defparam prom_inst_1.INIT_RAM_14 = 256'h5454545454545454545454545454545454545454545454545454545454545454;
defparam prom_inst_1.INIT_RAM_15 = 256'h545454545454545454545450657F7F7F7F7F7F7F7F7F61505454545454545454;
defparam prom_inst_1.INIT_RAM_16 = 256'h5454545454545454545454545454545454545454545454545454545454545454;
defparam prom_inst_1.INIT_RAM_17 = 256'h5454545454545454545454544C617F7F7F7F7F7F7F7F61505454545454545454;
defparam prom_inst_1.INIT_RAM_18 = 256'h5454545454545454545454545454545454545454545454545454545454545454;
defparam prom_inst_1.INIT_RAM_19 = 256'h5454545454545454545454545450617F7F7F7F7F7F7F61505454545454545454;
defparam prom_inst_1.INIT_RAM_1A = 256'h5050505050505050505050505050545454545454545454545454545454545454;
defparam prom_inst_1.INIT_RAM_1B = 256'h54545454545454545454545454544C617F7F7F7F7F7F5D4C5050505050505050;
defparam prom_inst_1.INIT_RAM_1C = 256'h6565656565656565656565656561545454545454545454545454545454545454;
defparam prom_inst_1.INIT_RAM_1D = 256'h5454545454545454545454545454544C617F7F7F7F7F6A5D6565656565656565;
defparam prom_inst_1.INIT_RAM_1E = 256'h7F7F7F7F7F7F7F7F7F7F7F7F7F7F5D5054545454545454545454545454545454;
defparam prom_inst_1.INIT_RAM_1F = 256'h545454545454545454545454545454544C617F7F7F7F7F7F7F7F7F7F7F7F7F7F;
defparam prom_inst_1.INIT_RAM_20 = 256'h7F7F7F7F7F7F7F7F7F7F7F7F7F7F5C5054545454545454545454545454545454;
defparam prom_inst_1.INIT_RAM_21 = 256'h54545454545454545454545454545454544C617F7F7F7F7F7F7F7F7F7F7F7F7F;
defparam prom_inst_1.INIT_RAM_22 = 256'h7F7F7F7F7F7F7F7F7F7F7F7F7F7F5C5054545454545454545454545454545454;
defparam prom_inst_1.INIT_RAM_23 = 256'h5454545454545454545454545454545454544C617F7F7F7F7F7F7F7F7F7F7F7F;
defparam prom_inst_1.INIT_RAM_24 = 256'h7F7F7F7F7F7F7F7F7F7F7F7F7F7F5C5054545454545454545454545454545454;
defparam prom_inst_1.INIT_RAM_25 = 256'h545454545454545454545454545454545454544C617F7F7F7F7F7F7F7F7F7F7F;
defparam prom_inst_1.INIT_RAM_26 = 256'h7F7F7F7F7F7F7F7F7F7F7F7F7F7F5C5054545454545454545454545454545454;
defparam prom_inst_1.INIT_RAM_27 = 256'h54545454545454545454545454545454545454544C617F7F7F7F7F7F7F7F7F7F;
defparam prom_inst_1.INIT_RAM_28 = 256'h7F7F7F7F7F7F7F7F7F7F7F7F7F7F5C5054545454545454545454545454545454;
defparam prom_inst_1.INIT_RAM_29 = 256'h5454545454545454545454545454545454545454544C617F7F7F7F7F7F7F7F7F;
defparam prom_inst_1.INIT_RAM_2A = 256'h7F7F7F7F7F7F7F7F7F7F7F7F7F7F5C5054545454545454545454545454545454;
defparam prom_inst_1.INIT_RAM_2B = 256'h545454545454545454545454545454545454545454544C617F7F7F7F7F7F7F7F;
defparam prom_inst_1.INIT_RAM_2C = 256'h7F7F7F7F7F7F7F7F7F7F7F7F7F7F5D5054545454545454545454545454545454;
defparam prom_inst_1.INIT_RAM_2D = 256'h54545454545454545454545454545454545454545454544C617F7F7F7F7F7F7F;
defparam prom_inst_1.INIT_RAM_2E = 256'h6E6E6E6E6E6E6E6E6E6E6E6E6E72585054545454545454545454545454545454;
defparam prom_inst_1.INIT_RAM_2F = 256'h5454545454545454545454545454545454545454545454545061726E6E6E6E6E;
defparam prom_inst_1.INIT_RAM_30 = 256'h4C4C4C4C4C4C4C4C4C4C4C4C4C50505454545454545454545454545454545054;
defparam prom_inst_1.INIT_RAM_31 = 256'h54545454545454545454545454545454545454545454545454504C4C4C4C4C4C;
defparam prom_inst_1.INIT_RAM_32 = 256'h5454545454545454545454545454545454545454545454545454545454545454;
defparam prom_inst_1.INIT_RAM_33 = 256'h5454545454545454545454545454545454545454545454545454545454545454;
defparam prom_inst_1.INIT_RAM_34 = 256'h5454545454545454545454545454545454545454545454545454545454545454;
defparam prom_inst_1.INIT_RAM_35 = 256'h5054545454545454545454545454545454545454545454545454545454545454;
defparam prom_inst_1.INIT_RAM_36 = 256'h545454545454545454545454545454545454545454545454545454545454505D;
defparam prom_inst_1.INIT_RAM_37 = 256'h5454545454545454545454545454545454545454545454545454545454545454;
defparam prom_inst_1.INIT_RAM_38 = 256'h5454545454545454545454545454545454545454545454545454545454545073;
defparam prom_inst_1.INIT_RAM_39 = 256'h6A50545454545454545454545454545454545454545454545454545454545454;
defparam prom_inst_1.INIT_RAM_3A = 256'h54545454545454545454545454545454545454545454545454545454544C657F;
defparam prom_inst_1.INIT_RAM_3B = 256'h7F614C5454545454545454545454545454545454545454545454545454545454;
defparam prom_inst_1.INIT_RAM_3C = 256'h5454545454545454545454545454545454545454545454545454545050657F7F;
defparam prom_inst_1.INIT_RAM_3D = 256'h7F7F615050545454545454545454545454545454545454545454545454545454;
defparam prom_inst_1.INIT_RAM_3E = 256'h5454545454545454545454545454545454545454545454545454545D737F7F7F;
defparam prom_inst_1.INIT_RAM_3F = 256'h7F7F7F6E5D545454545454545454545454545454545454545454545454545454;

pROM prom_inst_2 (
    .DO({prom_inst_2_dout_w[23:0],dout[23:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_2.READ_MODE = 1'b0;
defparam prom_inst_2.BIT_WIDTH = 8;
defparam prom_inst_2.RESET_MODE = "SYNC";
defparam prom_inst_2.INIT_RAM_00 = 256'h000000000000000000000000000000000000000000000000000000C5B4BBBBBB;
defparam prom_inst_2.INIT_RAM_01 = 256'hBBBBBB5284000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_02 = 256'h00000000000000000000000000000000000000000000000000000000006CBBBB;
defparam prom_inst_2.INIT_RAM_03 = 256'hBBBB080000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000008CBB;
defparam prom_inst_2.INIT_RAM_05 = 256'hBB08000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_06 = 256'h00000000000000000000000000000000000000000000000000000000000000D6;
defparam prom_inst_2.INIT_RAM_07 = 256'h5100000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000029;
defparam prom_inst_2.INIT_RAM_09 = 256'hA400000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000041;
defparam prom_inst_2.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_0E = 256'h000000000000000000000000000000000000AC1659F549000000000000000000;
defparam prom_inst_2.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_10 = 256'h0000000000000000000000000000000000B3FEFEFEFEFE0F0000000000000000;
defparam prom_inst_2.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_12 = 256'h7272727272A400000000000000000000CDFEFC162F58FCFD0700000000000000;
defparam prom_inst_2.INIT_RAM_13 = 256'h000000000000000000000000000000006B947272727272727272727272727272;
defparam prom_inst_2.INIT_RAM_14 = 256'hFDFDFDFDFE9A8400000000000000000016FE1600006379FE7200000000000000;
defparam prom_inst_2.INIT_RAM_15 = 256'h0000000000000000000000000000000072FFFDFDFDFDFDFDFDFDFDFDFDFDFDFD;
defparam prom_inst_2.INIT_RAM_16 = 256'hBBBBBBBBBAFD9A84000000000000000059FE51000000F5FED400000000000000;
defparam prom_inst_2.INIT_RAM_17 = 256'h0000000000000000000000000000000030FDBBBBBBBBBBBBBBBBBBBBBBBBBBBB;
defparam prom_inst_2.INIT_RAM_18 = 256'hBBBBBBBBBBBAFD9A8400000000000000F5FE586300E6BBFE5000000000000000;
defparam prom_inst_2.INIT_RAM_19 = 256'h0000000000000000000000000000000030FDBBBBBBBBBBBBBBBBBBBBBBBBBBBB;
defparam prom_inst_2.INIT_RAM_1A = 256'hBBBBBBBBBBBBBAFD9A840000000000004AFEDC99F4BBFCFCC500000000000000;
defparam prom_inst_2.INIT_RAM_1B = 256'h0000000000000000000000000000000030FDBBBBBBBBBBBBBBBBBBBBBBBBBBBB;
defparam prom_inst_2.INIT_RAM_1C = 256'hBBBBBBBBBBBBBBBAFD9A840000000000002FFDFEFEFEFC8B0000000000000000;
defparam prom_inst_2.INIT_RAM_1D = 256'h0000000000000000000000000000000030FDBBBBBBBBBBBBBBBBBBBBBBBBBBBB;
defparam prom_inst_2.INIT_RAM_1E = 256'hBBBBBBBBBBBBBBBBBAFD9A840000000000000792D551C5000000000000000000;
defparam prom_inst_2.INIT_RAM_1F = 256'h0000000000000000000000000000000030FDBBBBBBBBBBBBBBBBBBBBBBBBBBBB;
defparam prom_inst_2.INIT_RAM_20 = 256'hBABABABABABABABABBBAFD9A8400000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_21 = 256'h0000000000000000000000000000000030FDBABABABABABABABABABABABABABA;
defparam prom_inst_2.INIT_RAM_22 = 256'hFDFDFDFDFDFDFDFDDBBABAFD9A84000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_23 = 256'h0000000000000000000000000000000072FFFDFDFDFDFDFDFDFDFDFDFDFDFDFD;
defparam prom_inst_2.INIT_RAM_24 = 256'hACACACACACACAC8B37DCBBBAFD9A840000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_25 = 256'h0000000000000000000000000000000007CDACACACACACACACACACACACACACAC;
defparam prom_inst_2.INIT_RAM_26 = 256'h0000000000000000B4FDBBBBBAFD9A8400000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_28 = 256'h0000000000000000B4FCBBBBBBBAFD9A84000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_2A = 256'h0000000000000000B4FDBBBBBBBBBAFD9A840000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_2C = 256'h0000000000000000B4FDBBBBBBBBBBBAFD9BC500000000000000000000000000;
defparam prom_inst_2.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_2E = 256'h0000000000000000B4FDBBBBBBBBBBBABBFFCC00000000000000000000000000;
defparam prom_inst_2.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_30 = 256'h0000000000000000B4FDBBBBBBBBBABBFDCD0000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_32 = 256'h0000000000000000B4FDBBBBBBBABBFECD000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_34 = 256'h0000000000000000B3FCBBBBBABBFDCD00000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_36 = 256'h4242424242424200D4FCBBBABBFECD0000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000424242424242;
defparam prom_inst_2.INIT_RAM_38 = 256'h9A9A9A9A9A9A9A79BBBBBABBFDCC000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000093BB9A9A9A9A9A;
defparam prom_inst_2.INIT_RAM_3A = 256'hDBDBDBDBDBDBDBDCBBBABBFECD00000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_3B = 256'h000000000000000000000000000000000000000000000000B2FDDBDBDBDBDBDB;
defparam prom_inst_2.INIT_RAM_3C = 256'hBBBBBBBBBBBBBBBBBABBFDCC0000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000B3FDBBBBBBBBBBBBBB;
defparam prom_inst_2.INIT_RAM_3E = 256'hBBBBBBBBBBBBBBBABBFECD000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_3F = 256'h00000000000000000000000000000000000000000000B3FDBBBBBBBBBBBBBBBB;

pROM prom_inst_3 (
    .DO({prom_inst_3_dout_w[23:0],dout[31:24]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_3.READ_MODE = 1'b0;
defparam prom_inst_3.BIT_WIDTH = 8;
defparam prom_inst_3.RESET_MODE = "SYNC";
defparam prom_inst_3.INIT_RAM_00 = 256'h545454545454545454545454545454545454545454545454545450586E7F7F7F;
defparam prom_inst_3.INIT_RAM_01 = 256'h7F7F7F6A54505454545454545454545454545454545454545454545454545454;
defparam prom_inst_3.INIT_RAM_02 = 256'h5454545454545454545454545454545454545454545454545454545050617F7F;
defparam prom_inst_3.INIT_RAM_03 = 256'h7F7F5D5050545454545454545454545454545454545454545454545454545454;
defparam prom_inst_3.INIT_RAM_04 = 256'h54545454545454545454545454545454545454545454545454545454544C617F;
defparam prom_inst_3.INIT_RAM_05 = 256'h7F594C5454545454545454545454545454545454545454545454545454545454;
defparam prom_inst_3.INIT_RAM_06 = 256'h545454545454545454545454545454545454545454545454545454545454506E;
defparam prom_inst_3.INIT_RAM_07 = 256'h6A4C545454545454545454545454545454545454545454545454545454545454;
defparam prom_inst_3.INIT_RAM_08 = 256'h545454545454545454545454545454545454545454545454545454545454505D;
defparam prom_inst_3.INIT_RAM_09 = 256'h5854545454545454545454545454545454545454545454545454545454545454;
defparam prom_inst_3.INIT_RAM_0A = 256'h5454545454545454545454545454545454545450545454545454545454545454;
defparam prom_inst_3.INIT_RAM_0B = 256'h5454545454545454545454545454545454545454545454545454545454545454;
defparam prom_inst_3.INIT_RAM_0C = 256'h5454545454545454545454545454545454505050505050545454545454545054;
defparam prom_inst_3.INIT_RAM_0D = 256'h5454545454545454545454545454545454545454545454545454545454545454;
defparam prom_inst_3.INIT_RAM_0E = 256'h54545454545454545454545454545454505061777B76614C5454545454545454;
defparam prom_inst_3.INIT_RAM_0F = 256'h5454545454545454545454545454545454545454545454545454545454545454;
defparam prom_inst_3.INIT_RAM_10 = 256'h50505050505054545454545454545454506E7F7F7F7F7F665054545454545454;
defparam prom_inst_3.INIT_RAM_11 = 256'h54545454545454545454545454545454504C5050505050505050505050505050;
defparam prom_inst_3.INIT_RAM_12 = 256'h6E6E6E6E6E545054545454545454544C617F7F776A7B7F7F5D50545454545454;
defparam prom_inst_3.INIT_RAM_13 = 256'h5454545454545454545454545454545065726E6E6E6E6E6E6E6E6E6E6E6E6E6E;
defparam prom_inst_3.INIT_RAM_14 = 256'h7F7F7F7F7F7B54505454545454545450777F77504C507B7F6E50545454545454;
defparam prom_inst_3.INIT_RAM_15 = 256'h545454545454545454545454545454506E7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F;
defparam prom_inst_3.INIT_RAM_16 = 256'h7F7F7F7F7F7F7B5450545454545450547B7F6A48544C727F6E4C545454545454;
defparam prom_inst_3.INIT_RAM_17 = 256'h545454545454545454545454545454506E7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F;
defparam prom_inst_3.INIT_RAM_18 = 256'h7F7F7F7F7F7F7F7B5450545454545450727F7B544C587F7F6A4C545454545454;
defparam prom_inst_3.INIT_RAM_19 = 256'h545454545454545454545454545454506E7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F;
defparam prom_inst_3.INIT_RAM_1A = 256'h7F7F7F7F7F7F7F7F7B545054545454505D7F7F7B767F7F7F5850545454545454;
defparam prom_inst_3.INIT_RAM_1B = 256'h545454545454545454545454545454506E7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F;
defparam prom_inst_3.INIT_RAM_1C = 256'h7F7F7F7F7F7F7F7F7F7B54505454545450667F7F7F7F7F614C54545454545454;
defparam prom_inst_3.INIT_RAM_1D = 256'h545454545454545454545454545454506E7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F;
defparam prom_inst_3.INIT_RAM_1E = 256'h7F7F7F7F7F7F7F7F7F7F7B54505454545450596E766A58505454545454545454;
defparam prom_inst_3.INIT_RAM_1F = 256'h545454545454545454545454545454506E7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F;
defparam prom_inst_3.INIT_RAM_20 = 256'h7F7F7F7F7F7F7F7F7F7F7F7B5450545454545050505050545454545454545454;
defparam prom_inst_3.INIT_RAM_21 = 256'h545454545454545454545454545454506E7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F;
defparam prom_inst_3.INIT_RAM_22 = 256'h7F7F7F7F7F7F7F7F7F7F7F7F7B54505454545454545454545454545454545454;
defparam prom_inst_3.INIT_RAM_23 = 256'h545454545454545454545454545454506E7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F;
defparam prom_inst_3.INIT_RAM_24 = 256'h6161616161616161777F7F7F7F7B545054545454545454545454545454545454;
defparam prom_inst_3.INIT_RAM_25 = 256'h545454545454545454545454545454545D616161616161616161616161616161;
defparam prom_inst_3.INIT_RAM_26 = 256'h5050505050505048727F7F7F7F7F7B5450545454545454545454545454545454;
defparam prom_inst_3.INIT_RAM_27 = 256'h5454545454545454545454545454545450505050505050505050505050505050;
defparam prom_inst_3.INIT_RAM_28 = 256'h5454545454545450727F7F7F7F7F7F7B54505454545454545454545454545454;
defparam prom_inst_3.INIT_RAM_29 = 256'h5454545454545454545454545454545454545454545454545454545454545454;
defparam prom_inst_3.INIT_RAM_2A = 256'h545454545454544C727F7F7F7F7F7F7F7B545054545454545454545454545454;
defparam prom_inst_3.INIT_RAM_2B = 256'h5454545454545454545454545454545454545454545454545454545454545454;
defparam prom_inst_3.INIT_RAM_2C = 256'h545454545454544C727F7F7F7F7F7F7F7F7B5850545454545454545454545454;
defparam prom_inst_3.INIT_RAM_2D = 256'h5454545454545454545454545454545454545454545454545454545454545454;
defparam prom_inst_3.INIT_RAM_2E = 256'h545454545454544C727F7F7F7F7F7F7F7F7F6150505454545454545454545454;
defparam prom_inst_3.INIT_RAM_2F = 256'h5454545454545454545454545454545454545454545454545454545454545454;
defparam prom_inst_3.INIT_RAM_30 = 256'h545454545454544C727F7F7F7F7F7F7F7F655054545454545454545454545454;
defparam prom_inst_3.INIT_RAM_31 = 256'h5454545454545454545454545454545454545454545454545454545454545454;
defparam prom_inst_3.INIT_RAM_32 = 256'h545454545454544C727F7F7F7F7F7F7F65505454545454545454545454545454;
defparam prom_inst_3.INIT_RAM_33 = 256'h5454545454545454545454545454545454545454545454545454545454545454;
defparam prom_inst_3.INIT_RAM_34 = 256'h505050505050504C727F7F7F7F7F7F6550545454545454545454545454545454;
defparam prom_inst_3.INIT_RAM_35 = 256'h5454545454545454545454545454545454545454545454545454505050505050;
defparam prom_inst_3.INIT_RAM_36 = 256'h5454545454545450727F7F7F7F7F655054545454545454545454545454545454;
defparam prom_inst_3.INIT_RAM_37 = 256'h5454545454545454545454545454545454545454545454545050545454545454;
defparam prom_inst_3.INIT_RAM_38 = 256'h7F7F7F7F7F7F7F7F7F7F7F7F7F65505454545454545454545454545454545454;
defparam prom_inst_3.INIT_RAM_39 = 256'h545454545454545454545454545454545454545454545450506E7F7F7F7F7F7F;
defparam prom_inst_3.INIT_RAM_3A = 256'h7F7F7F7F7F7F7F7F7F7F7F7F6550545454545454545454545454545454545454;
defparam prom_inst_3.INIT_RAM_3B = 256'h54545454545454545454545454545454545454545454504C6E7F7F7F7F7F7F7F;
defparam prom_inst_3.INIT_RAM_3C = 256'h7F7F7F7F7F7F7F7F7F7F7F655050545454545454545454545454545454545454;
defparam prom_inst_3.INIT_RAM_3D = 256'h54545454545454545454545454545454545454545450506E7F7F7F7F7F7F7F7F;
defparam prom_inst_3.INIT_RAM_3E = 256'h7F7F7F7F7F7F7F7F7F7F65505454545454545454545454545454545454545454;
defparam prom_inst_3.INIT_RAM_3F = 256'h5454545454545454545454545454545454545454504C6E7F7F7F7F7F7F7F7F7F;

endmodule //Gowin_pROM
